seipp1@linux1.gl.umbc.edu.27067:1487878281