seipp1@linux1.gl.umbc.edu.20204:1487878281